library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port (
        clock : in std_logic;
        address_in : in unsigned(6 downto 0);
        data_out : out unsigned(15 downto 0)
    );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(15 downto 0);

    -- NOP         -> "0000"
    -- LD A, I     -> "0001"
    -- MOV A, Rn   -> "0010"
    -- MOV Rn, A   -> "0011"
    -- CMPI A, I   -> "0100"
    -- ADD A, Rn   -> "0101"
    -- SUB A, Rn   -> "0110"
    -- ADDI A, I   -> "0111"
    -- JMP address -> "1000"

    -- BHI offset_address -> "1001"
    -- BLT offset_address -> "1010"

    -- LW A, [Rn] -> "1011"
    -- SW [Rn], A -> "1100"
    
    constant rom_content : mem := (
        0 => B"0001_000000000000",
        1 => B"0111_000000000001",
        2 => B"0011_000_000000000",
        3 => B"1100_000_000000000",
        4 => B"0100_000000100000",
        5 => B"1010_00000_1111100",

        -- Zera múltiplos de 2
        6 => B"0001_000000000010",
        7 => B"0111_000000000010",
        8 => B"0011_000_000000000",
        9 => B"0001_000000000000",
        10 => B"1100_000_000000000",
        11 => B"0010_000_000000000",
        12 => B"0100_000000100000",
        13 => B"1010_00000_1111010",

        -- Zera múltiplos de 3
        14 => B"0001_000000000011",
        15 => B"0111_000000000011",
        16 => B"0011_000_000000000",
        17 => B"0001_000000000000",
        18 => B"1100_000_000000000",
        19 => B"0010_000_000000000",
        20 => B"0100_000000100000",
        21 => B"1010_00000_1111010",

        -- Zera múltiplos de 5
        22 => B"0001_000000000101",
        23 => B"0111_000000000101",
        24 => B"0011_000_000000000",
        25 => B"0001_000000000000",
        26 => B"1100_000_000000000",
        27 => B"0010_000_000000000",
        28 => B"0100_000000100000",
        29 => B"1010_00000_1111010",

        -- Zera múltiplos de 7
        30 => B"0001_000000000111",
        31 => B"0111_000000000111",
        32 => B"0011_000_000000000",
        33 => B"0001_000000000000",
        34 => B"1100_000_000000000",
        35 => B"0010_000_000000000",
        36 => B"0100_000000100000",
        37 => B"1010_00000_1111010",

        -- Zera múltiplos de 11
        38 => B"0001_000000001011",
        39 => B"0111_000000001011",
        40 => B"0011_000_000000000",
        41 => B"0001_000000000000",
        42 => B"1100_000_000000000",
        43 => B"0010_000_000000000",
        44 => B"0100_000000100000",
        45 => B"1010_00000_1111010",

        -- Zera múltiplos de 13
        46 => B"0001_000000001101",
        47 => B"0111_000000001101",
        48 => B"0011_000_000000000",
        49 => B"0001_000000000000",
        50 => B"1100_000_000000000",
        51 => B"0010_000_000000000",
        52 => B"0100_000000100000",
        53 => B"1010_00000_1111010",

        -- Zera múltiplos de 17
        54 => B"0001_000000010001",
        55 => B"0111_000000010001",
        56 => B"0011_000_000000000",
        57 => B"0001_000000000000",
        58 => B"1100_000_000000000",
        59 => B"0010_000_000000000",
        60 => B"0100_000000100000",
        61 => B"1010_00000_1111010",

        62 => B"0001_000000000001",
        63 => B"0111_000000000001",
        64 => B"0011_000_000000000",
        65 => B"1011_000_000000000",
        66 => B"0100_000000000000",
        67 => B"1001_00000_0000101",
        68 => B"0010_000_000000000",
        69 => B"0100_000000100000",
        70 => B"1010_00000_1111001",
        71 => B"1000_00000_1000111",
        72 => B"0011_001_000000000",
        73 => B"1000_00000_1000100",

        others => (others => '0')
    );

    -- constant rom_content : mem := (
    --     0 => B"0001_000001100100",
    --     1 => B"0011_000_000000000",
    --     2 => B"0001_000000010100",
    --     3 => B"0011_001_000000000",
    --     4 => B"0010_000_000000000",
    --     5 => B"1100_001_000000000",
    --     6 => B"0001_000011001000",
    --     7 => B"0011_000_000000000",
    --     8 => B"0001_000000101000",
    --     9 => B"0011_010_000000000",
    --     10 => B"0010_000_000000000",
    --     11 => B"1100_010_000000000",
    --     12 => B"1011_001_000000000",
    --     13 => B"1011_010_000000000",
    --     14 => B"1000_00000_0001110",
    --     others => (others => '0')
    -- );

    -- constant rom_content : mem := (
    --     0 => B"0001_000000000000",
    --     1 => B"0011_010_000000000",
    --     2 => B"0011_011_000000000",
    --     3 => B"0010_010_000000000",
    --     4 => B"0101_011_000000000",
    --     5 => B"0011_011_000000000",
    --     6 => B"0010_010_000000000",
    --     7 => B"0111_000000000001",
    --     8 => B"0011_010_000000000",
    --     9 => B"0100_000000011110",
    --     10 => B"1010_00000_1111001",
    --     11 => B"0010_011_000000000",
    --     12 => B"0011_100_000000000",
    --     others => (others => '0')
    -- );

    -- constant rom_content : mem := (
    --     0 => B"0001_000000000101",
    --     1 => B"0011_010_000000000",
    --     2 => B"0111_000000000011",
    --     3 => B"0011_011_000000000",
    --     4 => B"0010_010_000000000",
    --     5 => B"0101_011_000000000",
    --     6 => B"0011_100_000000000",
    --     7 => B"0111_111111111111",
    --     8 => B"0011_100_000000000",
    --     9 => B"1000_00000_0010100",
    --     10 => B"0001_000000000000",
    --     11 => B"0011_100_000000000",
    --     12 => B"0000_000000000000",
    --     13 => B"0000_000000000000",
    --     14 => B"0000_000000000000",
    --     15 => B"0000_000000000000",
    --     16 => B"0000_000000000000",
    --     17 => B"0000_000000000000",
    --     18 => B"0000_000000000000",
    --     19 => B"0000_000000000000",
    --     20 => B"0010_100_000000000",
    --     21 => B"0011_010_000000000",
    --     22 => B"1000_00000_0000100",
    --     23 => B"0001_000000000000",
    --     24 => B"0011_010_000000000",
    --     others => (others => '0')
    -- );
begin
    process(clock)
    begin
        if (rising_edge(clock)) then
            data_out <= rom_content(to_integer(address_in));
        end if;
    end process;
end architecture;